// SR Flip Flop
module srff(s, r, clk, rst, q, qbar);
  input s, r, clk, rst;
  output reg q, qbar;
  always @(posedge clk)
    begin
      if(rst == 1)
        begin
          q = 0; qbar = 1;
        end
      else
        begin
          case ({s, r})
            2'b00 : begin q = q; qbar = ~q ; end
            2'b01 : begin q = 1'b0; qbar = 1'b1 ; end
            2'b10 : begin q = 1'b1; qbar = 1'b0 ; end
            2'b11 : begin q = 1'bx; qbar = 1'bx ; end
          endcase
        end
    end
endmodule
